library verilog;
use verilog.vl_types.all;
entity fin_vlg_vec_tst is
end fin_vlg_vec_tst;
